package types;
    typedef enum {ALU_OP_ADD, ALU_OP_LT, ALU_OP_BOOL, ALU_OP_SHIFT} alu_op_t;

    // typedef enum bit [1:0] {
    //     BOOL_OP_XOR = 2'b00,
    //     BOOL_OP_NOR = 2'b01,
    //     BOOL_OP_OR = 2'b10,
    //     BOOL_OP_AND = 2'b11
    // } bool_op_t;
endpackage
